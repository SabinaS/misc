../lab1/camtest.sv