../lab1/write.sv