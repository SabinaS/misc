../lab1/cam.sv