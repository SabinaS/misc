../lab1/search.sv