../lab1/eff.sv