module camtest();

reg[]
